// Verilog netlist created by TD v5.0.29524
// Wed Mar 30 15:37:48 2022

`timescale 1ns / 1ps
module img_cache  // img_cache.v(14)
  (
  addra,
  addrb,
  cea,
  ceb,
  clka,
  clkb,
  dia,
  dob
  );

  input [15:0] addra;  // img_cache.v(35)
  input [15:0] addrb;  // img_cache.v(36)
  input cea;  // img_cache.v(37)
  input ceb;  // img_cache.v(38)
  input clka;  // img_cache.v(39)
  input clkb;  // img_cache.v(40)
  input [15:0] dia;  // img_cache.v(34)
  output [15:0] dob;  // img_cache.v(31)

  parameter ADDR_WIDTH_A = 16;
  parameter ADDR_WIDTH_B = 16;
  parameter DATA_DEPTH_A = 32800;
  parameter DATA_DEPTH_B = 32800;
  parameter DATA_WIDTH_A = 16;
  parameter DATA_WIDTH_B = 16;
  parameter REGMODE_A = "NOREG";
  parameter REGMODE_B = "NOREG";
  parameter WRITEMODE_A = "NORMAL";
  parameter WRITEMODE_B = "NORMAL";
  wire [0:6] addrb_piped;
  wire  \inst_dob_mux_b0/B1_0 ;
  wire  \inst_dob_mux_b0/B1_1 ;
  wire  \inst_dob_mux_b0/B1_10 ;
  wire  \inst_dob_mux_b0/B1_11 ;
  wire  \inst_dob_mux_b0/B1_12 ;
  wire  \inst_dob_mux_b0/B1_13 ;
  wire  \inst_dob_mux_b0/B1_14 ;
  wire  \inst_dob_mux_b0/B1_15 ;
  wire  \inst_dob_mux_b0/B1_2 ;
  wire  \inst_dob_mux_b0/B1_3 ;
  wire  \inst_dob_mux_b0/B1_4 ;
  wire  \inst_dob_mux_b0/B1_5 ;
  wire  \inst_dob_mux_b0/B1_6 ;
  wire  \inst_dob_mux_b0/B1_7 ;
  wire  \inst_dob_mux_b0/B1_8 ;
  wire  \inst_dob_mux_b0/B1_9 ;
  wire  \inst_dob_mux_b0/B2_0 ;
  wire  \inst_dob_mux_b0/B2_1 ;
  wire  \inst_dob_mux_b0/B2_2 ;
  wire  \inst_dob_mux_b0/B2_3 ;
  wire  \inst_dob_mux_b0/B2_4 ;
  wire  \inst_dob_mux_b0/B2_5 ;
  wire  \inst_dob_mux_b0/B2_6 ;
  wire  \inst_dob_mux_b0/B2_7 ;
  wire  \inst_dob_mux_b0/B3_0 ;
  wire  \inst_dob_mux_b0/B3_1 ;
  wire  \inst_dob_mux_b0/B3_2 ;
  wire  \inst_dob_mux_b0/B3_3 ;
  wire  \inst_dob_mux_b0/B4_0 ;
  wire  \inst_dob_mux_b0/B4_1 ;
  wire  \inst_dob_mux_b0/B5_0 ;
  wire  \inst_dob_mux_b1/B1_0 ;
  wire  \inst_dob_mux_b1/B1_1 ;
  wire  \inst_dob_mux_b1/B1_10 ;
  wire  \inst_dob_mux_b1/B1_11 ;
  wire  \inst_dob_mux_b1/B1_12 ;
  wire  \inst_dob_mux_b1/B1_13 ;
  wire  \inst_dob_mux_b1/B1_14 ;
  wire  \inst_dob_mux_b1/B1_15 ;
  wire  \inst_dob_mux_b1/B1_2 ;
  wire  \inst_dob_mux_b1/B1_3 ;
  wire  \inst_dob_mux_b1/B1_4 ;
  wire  \inst_dob_mux_b1/B1_5 ;
  wire  \inst_dob_mux_b1/B1_6 ;
  wire  \inst_dob_mux_b1/B1_7 ;
  wire  \inst_dob_mux_b1/B1_8 ;
  wire  \inst_dob_mux_b1/B1_9 ;
  wire  \inst_dob_mux_b1/B2_0 ;
  wire  \inst_dob_mux_b1/B2_1 ;
  wire  \inst_dob_mux_b1/B2_2 ;
  wire  \inst_dob_mux_b1/B2_3 ;
  wire  \inst_dob_mux_b1/B2_4 ;
  wire  \inst_dob_mux_b1/B2_5 ;
  wire  \inst_dob_mux_b1/B2_6 ;
  wire  \inst_dob_mux_b1/B2_7 ;
  wire  \inst_dob_mux_b1/B3_0 ;
  wire  \inst_dob_mux_b1/B3_1 ;
  wire  \inst_dob_mux_b1/B3_2 ;
  wire  \inst_dob_mux_b1/B3_3 ;
  wire  \inst_dob_mux_b1/B4_0 ;
  wire  \inst_dob_mux_b1/B4_1 ;
  wire  \inst_dob_mux_b1/B5_0 ;
  wire  \inst_dob_mux_b10/B4_0 ;
  wire  \inst_dob_mux_b10/B4_1 ;
  wire  \inst_dob_mux_b10/B5_0 ;
  wire  \inst_dob_mux_b11/B4_0 ;
  wire  \inst_dob_mux_b11/B4_1 ;
  wire  \inst_dob_mux_b11/B5_0 ;
  wire  \inst_dob_mux_b12/B4_0 ;
  wire  \inst_dob_mux_b12/B4_1 ;
  wire  \inst_dob_mux_b12/B5_0 ;
  wire  \inst_dob_mux_b13/B4_0 ;
  wire  \inst_dob_mux_b13/B4_1 ;
  wire  \inst_dob_mux_b13/B5_0 ;
  wire  \inst_dob_mux_b14/B4_0 ;
  wire  \inst_dob_mux_b14/B4_1 ;
  wire  \inst_dob_mux_b14/B5_0 ;
  wire  \inst_dob_mux_b15/B4_0 ;
  wire  \inst_dob_mux_b15/B4_1 ;
  wire  \inst_dob_mux_b15/B5_0 ;
  wire  \inst_dob_mux_b2/B1_0 ;
  wire  \inst_dob_mux_b2/B1_1 ;
  wire  \inst_dob_mux_b2/B1_10 ;
  wire  \inst_dob_mux_b2/B1_11 ;
  wire  \inst_dob_mux_b2/B1_12 ;
  wire  \inst_dob_mux_b2/B1_13 ;
  wire  \inst_dob_mux_b2/B1_14 ;
  wire  \inst_dob_mux_b2/B1_15 ;
  wire  \inst_dob_mux_b2/B1_2 ;
  wire  \inst_dob_mux_b2/B1_3 ;
  wire  \inst_dob_mux_b2/B1_4 ;
  wire  \inst_dob_mux_b2/B1_5 ;
  wire  \inst_dob_mux_b2/B1_6 ;
  wire  \inst_dob_mux_b2/B1_7 ;
  wire  \inst_dob_mux_b2/B1_8 ;
  wire  \inst_dob_mux_b2/B1_9 ;
  wire  \inst_dob_mux_b2/B2_0 ;
  wire  \inst_dob_mux_b2/B2_1 ;
  wire  \inst_dob_mux_b2/B2_2 ;
  wire  \inst_dob_mux_b2/B2_3 ;
  wire  \inst_dob_mux_b2/B2_4 ;
  wire  \inst_dob_mux_b2/B2_5 ;
  wire  \inst_dob_mux_b2/B2_6 ;
  wire  \inst_dob_mux_b2/B2_7 ;
  wire  \inst_dob_mux_b2/B3_0 ;
  wire  \inst_dob_mux_b2/B3_1 ;
  wire  \inst_dob_mux_b2/B3_2 ;
  wire  \inst_dob_mux_b2/B3_3 ;
  wire  \inst_dob_mux_b2/B4_0 ;
  wire  \inst_dob_mux_b2/B4_1 ;
  wire  \inst_dob_mux_b2/B5_0 ;
  wire  \inst_dob_mux_b3/B1_0 ;
  wire  \inst_dob_mux_b3/B1_1 ;
  wire  \inst_dob_mux_b3/B1_10 ;
  wire  \inst_dob_mux_b3/B1_11 ;
  wire  \inst_dob_mux_b3/B1_12 ;
  wire  \inst_dob_mux_b3/B1_13 ;
  wire  \inst_dob_mux_b3/B1_14 ;
  wire  \inst_dob_mux_b3/B1_15 ;
  wire  \inst_dob_mux_b3/B1_2 ;
  wire  \inst_dob_mux_b3/B1_3 ;
  wire  \inst_dob_mux_b3/B1_4 ;
  wire  \inst_dob_mux_b3/B1_5 ;
  wire  \inst_dob_mux_b3/B1_6 ;
  wire  \inst_dob_mux_b3/B1_7 ;
  wire  \inst_dob_mux_b3/B1_8 ;
  wire  \inst_dob_mux_b3/B1_9 ;
  wire  \inst_dob_mux_b3/B2_0 ;
  wire  \inst_dob_mux_b3/B2_1 ;
  wire  \inst_dob_mux_b3/B2_2 ;
  wire  \inst_dob_mux_b3/B2_3 ;
  wire  \inst_dob_mux_b3/B2_4 ;
  wire  \inst_dob_mux_b3/B2_5 ;
  wire  \inst_dob_mux_b3/B2_6 ;
  wire  \inst_dob_mux_b3/B2_7 ;
  wire  \inst_dob_mux_b3/B3_0 ;
  wire  \inst_dob_mux_b3/B3_1 ;
  wire  \inst_dob_mux_b3/B3_2 ;
  wire  \inst_dob_mux_b3/B3_3 ;
  wire  \inst_dob_mux_b3/B4_0 ;
  wire  \inst_dob_mux_b3/B4_1 ;
  wire  \inst_dob_mux_b3/B5_0 ;
  wire  \inst_dob_mux_b4/B1_0 ;
  wire  \inst_dob_mux_b4/B1_1 ;
  wire  \inst_dob_mux_b4/B1_10 ;
  wire  \inst_dob_mux_b4/B1_11 ;
  wire  \inst_dob_mux_b4/B1_12 ;
  wire  \inst_dob_mux_b4/B1_13 ;
  wire  \inst_dob_mux_b4/B1_14 ;
  wire  \inst_dob_mux_b4/B1_15 ;
  wire  \inst_dob_mux_b4/B1_2 ;
  wire  \inst_dob_mux_b4/B1_3 ;
  wire  \inst_dob_mux_b4/B1_4 ;
  wire  \inst_dob_mux_b4/B1_5 ;
  wire  \inst_dob_mux_b4/B1_6 ;
  wire  \inst_dob_mux_b4/B1_7 ;
  wire  \inst_dob_mux_b4/B1_8 ;
  wire  \inst_dob_mux_b4/B1_9 ;
  wire  \inst_dob_mux_b4/B2_0 ;
  wire  \inst_dob_mux_b4/B2_1 ;
  wire  \inst_dob_mux_b4/B2_2 ;
  wire  \inst_dob_mux_b4/B2_3 ;
  wire  \inst_dob_mux_b4/B2_4 ;
  wire  \inst_dob_mux_b4/B2_5 ;
  wire  \inst_dob_mux_b4/B2_6 ;
  wire  \inst_dob_mux_b4/B2_7 ;
  wire  \inst_dob_mux_b4/B3_0 ;
  wire  \inst_dob_mux_b4/B3_1 ;
  wire  \inst_dob_mux_b4/B3_2 ;
  wire  \inst_dob_mux_b4/B3_3 ;
  wire  \inst_dob_mux_b4/B4_0 ;
  wire  \inst_dob_mux_b4/B4_1 ;
  wire  \inst_dob_mux_b4/B5_0 ;
  wire  \inst_dob_mux_b5/B1_0 ;
  wire  \inst_dob_mux_b5/B1_1 ;
  wire  \inst_dob_mux_b5/B1_10 ;
  wire  \inst_dob_mux_b5/B1_11 ;
  wire  \inst_dob_mux_b5/B1_12 ;
  wire  \inst_dob_mux_b5/B1_13 ;
  wire  \inst_dob_mux_b5/B1_14 ;
  wire  \inst_dob_mux_b5/B1_15 ;
  wire  \inst_dob_mux_b5/B1_2 ;
  wire  \inst_dob_mux_b5/B1_3 ;
  wire  \inst_dob_mux_b5/B1_4 ;
  wire  \inst_dob_mux_b5/B1_5 ;
  wire  \inst_dob_mux_b5/B1_6 ;
  wire  \inst_dob_mux_b5/B1_7 ;
  wire  \inst_dob_mux_b5/B1_8 ;
  wire  \inst_dob_mux_b5/B1_9 ;
  wire  \inst_dob_mux_b5/B2_0 ;
  wire  \inst_dob_mux_b5/B2_1 ;
  wire  \inst_dob_mux_b5/B2_2 ;
  wire  \inst_dob_mux_b5/B2_3 ;
  wire  \inst_dob_mux_b5/B2_4 ;
  wire  \inst_dob_mux_b5/B2_5 ;
  wire  \inst_dob_mux_b5/B2_6 ;
  wire  \inst_dob_mux_b5/B2_7 ;
  wire  \inst_dob_mux_b5/B3_0 ;
  wire  \inst_dob_mux_b5/B3_1 ;
  wire  \inst_dob_mux_b5/B3_2 ;
  wire  \inst_dob_mux_b5/B3_3 ;
  wire  \inst_dob_mux_b5/B4_0 ;
  wire  \inst_dob_mux_b5/B4_1 ;
  wire  \inst_dob_mux_b5/B5_0 ;
  wire  \inst_dob_mux_b6/B1_0 ;
  wire  \inst_dob_mux_b6/B1_1 ;
  wire  \inst_dob_mux_b6/B1_10 ;
  wire  \inst_dob_mux_b6/B1_11 ;
  wire  \inst_dob_mux_b6/B1_12 ;
  wire  \inst_dob_mux_b6/B1_13 ;
  wire  \inst_dob_mux_b6/B1_14 ;
  wire  \inst_dob_mux_b6/B1_15 ;
  wire  \inst_dob_mux_b6/B1_2 ;
  wire  \inst_dob_mux_b6/B1_3 ;
  wire  \inst_dob_mux_b6/B1_4 ;
  wire  \inst_dob_mux_b6/B1_5 ;
  wire  \inst_dob_mux_b6/B1_6 ;
  wire  \inst_dob_mux_b6/B1_7 ;
  wire  \inst_dob_mux_b6/B1_8 ;
  wire  \inst_dob_mux_b6/B1_9 ;
  wire  \inst_dob_mux_b6/B2_0 ;
  wire  \inst_dob_mux_b6/B2_1 ;
  wire  \inst_dob_mux_b6/B2_2 ;
  wire  \inst_dob_mux_b6/B2_3 ;
  wire  \inst_dob_mux_b6/B2_4 ;
  wire  \inst_dob_mux_b6/B2_5 ;
  wire  \inst_dob_mux_b6/B2_6 ;
  wire  \inst_dob_mux_b6/B2_7 ;
  wire  \inst_dob_mux_b6/B3_0 ;
  wire  \inst_dob_mux_b6/B3_1 ;
  wire  \inst_dob_mux_b6/B3_2 ;
  wire  \inst_dob_mux_b6/B3_3 ;
  wire  \inst_dob_mux_b6/B4_0 ;
  wire  \inst_dob_mux_b6/B4_1 ;
  wire  \inst_dob_mux_b6/B5_0 ;
  wire  \inst_dob_mux_b7/B1_0 ;
  wire  \inst_dob_mux_b7/B1_1 ;
  wire  \inst_dob_mux_b7/B1_10 ;
  wire  \inst_dob_mux_b7/B1_11 ;
  wire  \inst_dob_mux_b7/B1_12 ;
  wire  \inst_dob_mux_b7/B1_13 ;
  wire  \inst_dob_mux_b7/B1_14 ;
  wire  \inst_dob_mux_b7/B1_15 ;
  wire  \inst_dob_mux_b7/B1_2 ;
  wire  \inst_dob_mux_b7/B1_3 ;
  wire  \inst_dob_mux_b7/B1_4 ;
  wire  \inst_dob_mux_b7/B1_5 ;
  wire  \inst_dob_mux_b7/B1_6 ;
  wire  \inst_dob_mux_b7/B1_7 ;
  wire  \inst_dob_mux_b7/B1_8 ;
  wire  \inst_dob_mux_b7/B1_9 ;
  wire  \inst_dob_mux_b7/B2_0 ;
  wire  \inst_dob_mux_b7/B2_1 ;
  wire  \inst_dob_mux_b7/B2_2 ;
  wire  \inst_dob_mux_b7/B2_3 ;
  wire  \inst_dob_mux_b7/B2_4 ;
  wire  \inst_dob_mux_b7/B2_5 ;
  wire  \inst_dob_mux_b7/B2_6 ;
  wire  \inst_dob_mux_b7/B2_7 ;
  wire  \inst_dob_mux_b7/B3_0 ;
  wire  \inst_dob_mux_b7/B3_1 ;
  wire  \inst_dob_mux_b7/B3_2 ;
  wire  \inst_dob_mux_b7/B3_3 ;
  wire  \inst_dob_mux_b7/B4_0 ;
  wire  \inst_dob_mux_b7/B4_1 ;
  wire  \inst_dob_mux_b7/B5_0 ;
  wire  \inst_dob_mux_b8/B1_0 ;
  wire  \inst_dob_mux_b8/B1_1 ;
  wire  \inst_dob_mux_b8/B1_10 ;
  wire  \inst_dob_mux_b8/B1_11 ;
  wire  \inst_dob_mux_b8/B1_12 ;
  wire  \inst_dob_mux_b8/B1_13 ;
  wire  \inst_dob_mux_b8/B1_14 ;
  wire  \inst_dob_mux_b8/B1_15 ;
  wire  \inst_dob_mux_b8/B1_2 ;
  wire  \inst_dob_mux_b8/B1_3 ;
  wire  \inst_dob_mux_b8/B1_4 ;
  wire  \inst_dob_mux_b8/B1_5 ;
  wire  \inst_dob_mux_b8/B1_6 ;
  wire  \inst_dob_mux_b8/B1_7 ;
  wire  \inst_dob_mux_b8/B1_8 ;
  wire  \inst_dob_mux_b8/B1_9 ;
  wire  \inst_dob_mux_b8/B2_0 ;
  wire  \inst_dob_mux_b8/B2_1 ;
  wire  \inst_dob_mux_b8/B2_2 ;
  wire  \inst_dob_mux_b8/B2_3 ;
  wire  \inst_dob_mux_b8/B2_4 ;
  wire  \inst_dob_mux_b8/B2_5 ;
  wire  \inst_dob_mux_b8/B2_6 ;
  wire  \inst_dob_mux_b8/B2_7 ;
  wire  \inst_dob_mux_b8/B3_0 ;
  wire  \inst_dob_mux_b8/B3_1 ;
  wire  \inst_dob_mux_b8/B3_2 ;
  wire  \inst_dob_mux_b8/B3_3 ;
  wire  \inst_dob_mux_b8/B4_0 ;
  wire  \inst_dob_mux_b8/B4_1 ;
  wire  \inst_dob_mux_b8/B5_0 ;
  wire  \inst_dob_mux_b9/B4_0 ;
  wire  \inst_dob_mux_b9/B4_1 ;
  wire  \inst_dob_mux_b9/B5_0 ;
  wire \and_Naddra[11]_Naddr_o ;
  wire \and_Naddra[11]_Naddr_o_and_cea ;
  wire \and_Naddra[12]_Naddr_o ;
  wire \and_Naddra[12]_Naddr_o_al_n54 ;
  wire \and_Naddra[12]_addra_o ;
  wire \and_Naddra[12]_addra_o_al_n86 ;
  wire \and_Naddrb[11]_Naddr_o ;
  wire \and_Naddrb[11]_Naddr_o_and_ceb ;
  wire \and_Naddrb[12]_Naddr_o ;
  wire \and_Naddrb[12]_Naddr_o_al_n57 ;
  wire \and_Naddrb[12]_addrb_o ;
  wire \and_Naddrb[12]_addrb_o_al_n89 ;
  wire \and_addra[12]_Naddra_o ;
  wire \and_addra[12]_Naddra_o_al_n70 ;
  wire \and_addra[12]_addra[_o ;
  wire \and_addra[12]_addra[_o_al_n102 ;
  wire \and_addrb[12]_Naddrb_o ;
  wire \and_addrb[12]_Naddrb_o_al_n73 ;
  wire \and_addrb[12]_addrb[_o ;
  wire \and_addrb[12]_addrb[_o_al_n105 ;
  wire inst_dob_i0_000;
  wire inst_dob_i0_001;
  wire inst_dob_i0_002;
  wire inst_dob_i0_003;
  wire inst_dob_i0_004;
  wire inst_dob_i0_005;
  wire inst_dob_i0_006;
  wire inst_dob_i0_007;
  wire inst_dob_i0_008;
  wire inst_dob_i0_009;
  wire inst_dob_i0_010;
  wire inst_dob_i0_011;
  wire inst_dob_i0_012;
  wire inst_dob_i0_013;
  wire inst_dob_i0_014;
  wire inst_dob_i0_015;
  wire inst_dob_i10_000;
  wire inst_dob_i10_001;
  wire inst_dob_i10_002;
  wire inst_dob_i10_003;
  wire inst_dob_i10_004;
  wire inst_dob_i10_005;
  wire inst_dob_i10_006;
  wire inst_dob_i10_007;
  wire inst_dob_i10_008;
  wire inst_dob_i12_000;
  wire inst_dob_i12_001;
  wire inst_dob_i12_002;
  wire inst_dob_i12_003;
  wire inst_dob_i12_004;
  wire inst_dob_i12_005;
  wire inst_dob_i12_006;
  wire inst_dob_i12_007;
  wire inst_dob_i12_008;
  wire inst_dob_i14_000;
  wire inst_dob_i14_001;
  wire inst_dob_i14_002;
  wire inst_dob_i14_003;
  wire inst_dob_i14_004;
  wire inst_dob_i14_005;
  wire inst_dob_i14_006;
  wire inst_dob_i14_007;
  wire inst_dob_i14_008;
  wire inst_dob_i16_000;
  wire inst_dob_i16_001;
  wire inst_dob_i16_002;
  wire inst_dob_i16_003;
  wire inst_dob_i16_004;
  wire inst_dob_i16_005;
  wire inst_dob_i16_006;
  wire inst_dob_i16_007;
  wire inst_dob_i16_008;
  wire inst_dob_i16_009;
  wire inst_dob_i16_010;
  wire inst_dob_i16_011;
  wire inst_dob_i16_012;
  wire inst_dob_i16_013;
  wire inst_dob_i16_014;
  wire inst_dob_i16_015;
  wire inst_dob_i18_000;
  wire inst_dob_i18_001;
  wire inst_dob_i18_002;
  wire inst_dob_i18_003;
  wire inst_dob_i18_004;
  wire inst_dob_i18_005;
  wire inst_dob_i18_006;
  wire inst_dob_i18_007;
  wire inst_dob_i18_008;
  wire inst_dob_i20_000;
  wire inst_dob_i20_001;
  wire inst_dob_i20_002;
  wire inst_dob_i20_003;
  wire inst_dob_i20_004;
  wire inst_dob_i20_005;
  wire inst_dob_i20_006;
  wire inst_dob_i20_007;
  wire inst_dob_i20_008;
  wire inst_dob_i22_000;
  wire inst_dob_i22_001;
  wire inst_dob_i22_002;
  wire inst_dob_i22_003;
  wire inst_dob_i22_004;
  wire inst_dob_i22_005;
  wire inst_dob_i22_006;
  wire inst_dob_i22_007;
  wire inst_dob_i22_008;
  wire inst_dob_i24_000;
  wire inst_dob_i24_001;
  wire inst_dob_i24_002;
  wire inst_dob_i24_003;
  wire inst_dob_i24_004;
  wire inst_dob_i24_005;
  wire inst_dob_i24_006;
  wire inst_dob_i24_007;
  wire inst_dob_i24_008;
  wire inst_dob_i26_000;
  wire inst_dob_i26_001;
  wire inst_dob_i26_002;
  wire inst_dob_i26_003;
  wire inst_dob_i26_004;
  wire inst_dob_i26_005;
  wire inst_dob_i26_006;
  wire inst_dob_i26_007;
  wire inst_dob_i26_008;
  wire inst_dob_i28_000;
  wire inst_dob_i28_001;
  wire inst_dob_i28_002;
  wire inst_dob_i28_003;
  wire inst_dob_i28_004;
  wire inst_dob_i28_005;
  wire inst_dob_i28_006;
  wire inst_dob_i28_007;
  wire inst_dob_i28_008;
  wire inst_dob_i2_000;
  wire inst_dob_i2_001;
  wire inst_dob_i2_002;
  wire inst_dob_i2_003;
  wire inst_dob_i2_004;
  wire inst_dob_i2_005;
  wire inst_dob_i2_006;
  wire inst_dob_i2_007;
  wire inst_dob_i2_008;
  wire inst_dob_i30_000;
  wire inst_dob_i30_001;
  wire inst_dob_i30_002;
  wire inst_dob_i30_003;
  wire inst_dob_i30_004;
  wire inst_dob_i30_005;
  wire inst_dob_i30_006;
  wire inst_dob_i30_007;
  wire inst_dob_i30_008;
  wire inst_dob_i32_000;
  wire inst_dob_i32_001;
  wire inst_dob_i32_002;
  wire inst_dob_i32_003;
  wire inst_dob_i32_004;
  wire inst_dob_i32_005;
  wire inst_dob_i32_006;
  wire inst_dob_i32_007;
  wire inst_dob_i32_008;
  wire inst_dob_i32_009;
  wire inst_dob_i32_010;
  wire inst_dob_i32_011;
  wire inst_dob_i32_012;
  wire inst_dob_i32_013;
  wire inst_dob_i32_014;
  wire inst_dob_i32_015;
  wire inst_dob_i34_000;
  wire inst_dob_i34_001;
  wire inst_dob_i34_002;
  wire inst_dob_i34_003;
  wire inst_dob_i34_004;
  wire inst_dob_i34_005;
  wire inst_dob_i34_006;
  wire inst_dob_i34_007;
  wire inst_dob_i34_008;
  wire inst_dob_i36_000;
  wire inst_dob_i36_001;
  wire inst_dob_i36_002;
  wire inst_dob_i36_003;
  wire inst_dob_i36_004;
  wire inst_dob_i36_005;
  wire inst_dob_i36_006;
  wire inst_dob_i36_007;
  wire inst_dob_i36_008;
  wire inst_dob_i38_000;
  wire inst_dob_i38_001;
  wire inst_dob_i38_002;
  wire inst_dob_i38_003;
  wire inst_dob_i38_004;
  wire inst_dob_i38_005;
  wire inst_dob_i38_006;
  wire inst_dob_i38_007;
  wire inst_dob_i38_008;
  wire inst_dob_i40_000;
  wire inst_dob_i40_001;
  wire inst_dob_i40_002;
  wire inst_dob_i40_003;
  wire inst_dob_i40_004;
  wire inst_dob_i40_005;
  wire inst_dob_i40_006;
  wire inst_dob_i40_007;
  wire inst_dob_i40_008;
  wire inst_dob_i42_000;
  wire inst_dob_i42_001;
  wire inst_dob_i42_002;
  wire inst_dob_i42_003;
  wire inst_dob_i42_004;
  wire inst_dob_i42_005;
  wire inst_dob_i42_006;
  wire inst_dob_i42_007;
  wire inst_dob_i42_008;
  wire inst_dob_i44_000;
  wire inst_dob_i44_001;
  wire inst_dob_i44_002;
  wire inst_dob_i44_003;
  wire inst_dob_i44_004;
  wire inst_dob_i44_005;
  wire inst_dob_i44_006;
  wire inst_dob_i44_007;
  wire inst_dob_i44_008;
  wire inst_dob_i46_000;
  wire inst_dob_i46_001;
  wire inst_dob_i46_002;
  wire inst_dob_i46_003;
  wire inst_dob_i46_004;
  wire inst_dob_i46_005;
  wire inst_dob_i46_006;
  wire inst_dob_i46_007;
  wire inst_dob_i46_008;
  wire inst_dob_i48_000;
  wire inst_dob_i48_001;
  wire inst_dob_i48_002;
  wire inst_dob_i48_003;
  wire inst_dob_i48_004;
  wire inst_dob_i48_005;
  wire inst_dob_i48_006;
  wire inst_dob_i48_007;
  wire inst_dob_i48_008;
  wire inst_dob_i48_009;
  wire inst_dob_i48_010;
  wire inst_dob_i48_011;
  wire inst_dob_i48_012;
  wire inst_dob_i48_013;
  wire inst_dob_i48_014;
  wire inst_dob_i48_015;
  wire inst_dob_i4_000;
  wire inst_dob_i4_001;
  wire inst_dob_i4_002;
  wire inst_dob_i4_003;
  wire inst_dob_i4_004;
  wire inst_dob_i4_005;
  wire inst_dob_i4_006;
  wire inst_dob_i4_007;
  wire inst_dob_i4_008;
  wire inst_dob_i50_000;
  wire inst_dob_i50_001;
  wire inst_dob_i50_002;
  wire inst_dob_i50_003;
  wire inst_dob_i50_004;
  wire inst_dob_i50_005;
  wire inst_dob_i50_006;
  wire inst_dob_i50_007;
  wire inst_dob_i50_008;
  wire inst_dob_i52_000;
  wire inst_dob_i52_001;
  wire inst_dob_i52_002;
  wire inst_dob_i52_003;
  wire inst_dob_i52_004;
  wire inst_dob_i52_005;
  wire inst_dob_i52_006;
  wire inst_dob_i52_007;
  wire inst_dob_i52_008;
  wire inst_dob_i54_000;
  wire inst_dob_i54_001;
  wire inst_dob_i54_002;
  wire inst_dob_i54_003;
  wire inst_dob_i54_004;
  wire inst_dob_i54_005;
  wire inst_dob_i54_006;
  wire inst_dob_i54_007;
  wire inst_dob_i54_008;
  wire inst_dob_i56_000;
  wire inst_dob_i56_001;
  wire inst_dob_i56_002;
  wire inst_dob_i56_003;
  wire inst_dob_i56_004;
  wire inst_dob_i56_005;
  wire inst_dob_i56_006;
  wire inst_dob_i56_007;
  wire inst_dob_i56_008;
  wire inst_dob_i58_000;
  wire inst_dob_i58_001;
  wire inst_dob_i58_002;
  wire inst_dob_i58_003;
  wire inst_dob_i58_004;
  wire inst_dob_i58_005;
  wire inst_dob_i58_006;
  wire inst_dob_i58_007;
  wire inst_dob_i58_008;
  wire inst_dob_i60_000;
  wire inst_dob_i60_001;
  wire inst_dob_i60_002;
  wire inst_dob_i60_003;
  wire inst_dob_i60_004;
  wire inst_dob_i60_005;
  wire inst_dob_i60_006;
  wire inst_dob_i60_007;
  wire inst_dob_i60_008;
  wire inst_dob_i62_000;
  wire inst_dob_i62_001;
  wire inst_dob_i62_002;
  wire inst_dob_i62_003;
  wire inst_dob_i62_004;
  wire inst_dob_i62_005;
  wire inst_dob_i62_006;
  wire inst_dob_i62_007;
  wire inst_dob_i62_008;
  wire inst_dob_i64_000;
  wire inst_dob_i64_001;
  wire inst_dob_i64_002;
  wire inst_dob_i64_003;
  wire inst_dob_i64_004;
  wire inst_dob_i64_005;
  wire inst_dob_i64_006;
  wire inst_dob_i64_007;
  wire inst_dob_i64_008;
  wire inst_dob_i64_009;
  wire inst_dob_i64_010;
  wire inst_dob_i64_011;
  wire inst_dob_i64_012;
  wire inst_dob_i64_013;
  wire inst_dob_i64_014;
  wire inst_dob_i64_015;
  wire inst_dob_i6_000;
  wire inst_dob_i6_001;
  wire inst_dob_i6_002;
  wire inst_dob_i6_003;
  wire inst_dob_i6_004;
  wire inst_dob_i6_005;
  wire inst_dob_i6_006;
  wire inst_dob_i6_007;
  wire inst_dob_i6_008;
  wire inst_dob_i8_000;
  wire inst_dob_i8_001;
  wire inst_dob_i8_002;
  wire inst_dob_i8_003;
  wire inst_dob_i8_004;
  wire inst_dob_i8_005;
  wire inst_dob_i8_006;
  wire inst_dob_i8_007;
  wire inst_dob_i8_008;

  AL_DFF_X addrb_pipe_b1 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[10]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[1]));
  AL_DFF_X addrb_pipe_b2 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[11]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[2]));
  AL_DFF_X addrb_pipe_b3 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[12]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[3]));
  AL_DFF_X addrb_pipe_b4 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[13]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[4]));
  AL_DFF_X addrb_pipe_b5 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[14]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[5]));
  AL_DFF_X addrb_pipe_b6 (
    .ar(1'b0),
    .as(1'b0),
    .clk(clkb),
    .d(addrb[15]),
    .en(ceb),
    .sr(1'b0),
    .ss(1'b0),
    .q(addrb_piped[6]));
  and \and_Naddra[11]_Naddr  (\and_Naddra[11]_Naddr_o , ~addra[11], ~addra[12], ~addra[13], ~addra[14], addra[15]);
  and \and_Naddra[11]_Naddr_o_and_cea_i  (\and_Naddra[11]_Naddr_o_and_cea , \and_Naddra[11]_Naddr_o , cea);
  and \and_Naddra[12]_Naddr  (\and_Naddra[12]_Naddr_o , ~addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_Naddr_al_u54  (\and_Naddra[12]_Naddr_o_al_n54 , ~addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_Naddra[12]_addra  (\and_Naddra[12]_addra_o , ~addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_Naddra[12]_addra_al_u86  (\and_Naddra[12]_addra_o_al_n86 , ~addra[12], addra[13], addra[14], ~addra[15]);
  and \and_Naddrb[11]_Naddr  (\and_Naddrb[11]_Naddr_o , ~addrb[11], ~addrb[12], ~addrb[13], ~addrb[14], addrb[15]);
  and \and_Naddrb[11]_Naddr_o_and_ceb_i  (\and_Naddrb[11]_Naddr_o_and_ceb , \and_Naddrb[11]_Naddr_o , ceb);
  and \and_Naddrb[12]_Naddr  (\and_Naddrb[12]_Naddr_o , ~addrb[12], ~addrb[13], ~addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_Naddr_al_u57  (\and_Naddrb[12]_Naddr_o_al_n57 , ~addrb[12], ~addrb[13], addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_addrb  (\and_Naddrb[12]_addrb_o , ~addrb[12], addrb[13], ~addrb[14], ~addrb[15]);
  and \and_Naddrb[12]_addrb_al_u89  (\and_Naddrb[12]_addrb_o_al_n89 , ~addrb[12], addrb[13], addrb[14], ~addrb[15]);
  and \and_addra[12]_Naddra  (\and_addra[12]_Naddra_o , addra[12], ~addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_Naddra_al_u70  (\and_addra[12]_Naddra_o_al_n70 , addra[12], ~addra[13], addra[14], ~addra[15]);
  and \and_addra[12]_addra[  (\and_addra[12]_addra[_o , addra[12], addra[13], ~addra[14], ~addra[15]);
  and \and_addra[12]_addra[_al_u102  (\and_addra[12]_addra[_o_al_n102 , addra[12], addra[13], addra[14], ~addra[15]);
  and \and_addrb[12]_Naddrb  (\and_addrb[12]_Naddrb_o , addrb[12], ~addrb[13], ~addrb[14], ~addrb[15]);
  and \and_addrb[12]_Naddrb_al_u73  (\and_addrb[12]_Naddrb_o_al_n73 , addrb[12], ~addrb[13], addrb[14], ~addrb[15]);
  and \and_addrb[12]_addrb[  (\and_addrb[12]_addrb[_o , addrb[12], addrb[13], ~addrb[14], ~addrb[15]);
  and \and_addrb[12]_addrb[_al_u105  (\and_addrb[12]_addrb[_o_al_n105 , addrb[12], addrb[13], addrb[14], ~addrb[15]);
  EG_PHY_CONFIG #(
    .DONE_PERSISTN("ENABLE"),
    .INIT_PERSISTN("ENABLE"),
    .JTAG_PERSISTN("DISABLE"),
    .PROGRAMN_PERSISTN("DISABLE"))
    config_inst ();
  // address_offset=0;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i0_008,inst_dob_i0_007,inst_dob_i0_006,inst_dob_i0_005,inst_dob_i0_004,inst_dob_i0_003,inst_dob_i0_002,inst_dob_i0_001,inst_dob_i0_000}));
  // address_offset=0;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n71,open_n72,open_n73,open_n74,open_n75,open_n76,open_n77,dia[9],open_n78}),
    .dob({open_n103,open_n104,open_n105,open_n106,open_n107,open_n108,open_n109,open_n110,inst_dob_i0_009}));
  // address_offset=0;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n111,open_n112,open_n113,open_n114,open_n115,open_n116,open_n117,dia[10],open_n118}),
    .dob({open_n143,open_n144,open_n145,open_n146,open_n147,open_n148,open_n149,open_n150,inst_dob_i0_010}));
  // address_offset=0;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n151,open_n152,open_n153,open_n154,open_n155,open_n156,open_n157,dia[11],open_n158}),
    .dob({open_n183,open_n184,open_n185,open_n186,open_n187,open_n188,open_n189,open_n190,inst_dob_i0_011}));
  // address_offset=0;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n191,open_n192,open_n193,open_n194,open_n195,open_n196,open_n197,dia[12],open_n198}),
    .dob({open_n223,open_n224,open_n225,open_n226,open_n227,open_n228,open_n229,open_n230,inst_dob_i0_012}));
  // address_offset=0;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n231,open_n232,open_n233,open_n234,open_n235,open_n236,open_n237,dia[13],open_n238}),
    .dob({open_n263,open_n264,open_n265,open_n266,open_n267,open_n268,open_n269,open_n270,inst_dob_i0_013}));
  // address_offset=0;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n271,open_n272,open_n273,open_n274,open_n275,open_n276,open_n277,dia[14],open_n278}),
    .dob({open_n303,open_n304,open_n305,open_n306,open_n307,open_n308,open_n309,open_n310,inst_dob_i0_014}));
  // address_offset=0;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_000000_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n311,open_n312,open_n313,open_n314,open_n315,open_n316,open_n317,dia[15],open_n318}),
    .dob({open_n343,open_n344,open_n345,open_n346,open_n347,open_n348,open_n349,open_n350,inst_dob_i0_015}));
  // address_offset=1024;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_001024_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i2_008,inst_dob_i2_007,inst_dob_i2_006,inst_dob_i2_005,inst_dob_i2_004,inst_dob_i2_003,inst_dob_i2_002,inst_dob_i2_001,inst_dob_i2_000}));
  // address_offset=2048;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_002048_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i4_008,inst_dob_i4_007,inst_dob_i4_006,inst_dob_i4_005,inst_dob_i4_004,inst_dob_i4_003,inst_dob_i4_002,inst_dob_i4_001,inst_dob_i4_000}));
  // address_offset=3072;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_003072_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i6_008,inst_dob_i6_007,inst_dob_i6_006,inst_dob_i6_005,inst_dob_i6_004,inst_dob_i6_003,inst_dob_i6_002,inst_dob_i6_001,inst_dob_i6_000}));
  // address_offset=4096;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_004096_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i8_008,inst_dob_i8_007,inst_dob_i8_006,inst_dob_i8_005,inst_dob_i8_004,inst_dob_i8_003,inst_dob_i8_002,inst_dob_i8_001,inst_dob_i8_000}));
  // address_offset=5120;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_005120_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i10_008,inst_dob_i10_007,inst_dob_i10_006,inst_dob_i10_005,inst_dob_i10_004,inst_dob_i10_003,inst_dob_i10_002,inst_dob_i10_001,inst_dob_i10_000}));
  // address_offset=6144;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_006144_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i12_008,inst_dob_i12_007,inst_dob_i12_006,inst_dob_i12_005,inst_dob_i12_004,inst_dob_i12_003,inst_dob_i12_002,inst_dob_i12_001,inst_dob_i12_000}));
  // address_offset=7168;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_007168_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i14_008,inst_dob_i14_007,inst_dob_i14_006,inst_dob_i14_005,inst_dob_i14_004,inst_dob_i14_003,inst_dob_i14_002,inst_dob_i14_001,inst_dob_i14_000}));
  // address_offset=8192;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i16_008,inst_dob_i16_007,inst_dob_i16_006,inst_dob_i16_005,inst_dob_i16_004,inst_dob_i16_003,inst_dob_i16_002,inst_dob_i16_001,inst_dob_i16_000}));
  // address_offset=8192;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n543,open_n544,open_n545,open_n546,open_n547,open_n548,open_n549,dia[9],open_n550}),
    .dob({open_n575,open_n576,open_n577,open_n578,open_n579,open_n580,open_n581,open_n582,inst_dob_i16_009}));
  // address_offset=8192;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n583,open_n584,open_n585,open_n586,open_n587,open_n588,open_n589,dia[10],open_n590}),
    .dob({open_n615,open_n616,open_n617,open_n618,open_n619,open_n620,open_n621,open_n622,inst_dob_i16_010}));
  // address_offset=8192;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n623,open_n624,open_n625,open_n626,open_n627,open_n628,open_n629,dia[11],open_n630}),
    .dob({open_n655,open_n656,open_n657,open_n658,open_n659,open_n660,open_n661,open_n662,inst_dob_i16_011}));
  // address_offset=8192;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n663,open_n664,open_n665,open_n666,open_n667,open_n668,open_n669,dia[12],open_n670}),
    .dob({open_n695,open_n696,open_n697,open_n698,open_n699,open_n700,open_n701,open_n702,inst_dob_i16_012}));
  // address_offset=8192;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n703,open_n704,open_n705,open_n706,open_n707,open_n708,open_n709,dia[13],open_n710}),
    .dob({open_n735,open_n736,open_n737,open_n738,open_n739,open_n740,open_n741,open_n742,inst_dob_i16_013}));
  // address_offset=8192;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n743,open_n744,open_n745,open_n746,open_n747,open_n748,open_n749,dia[14],open_n750}),
    .dob({open_n775,open_n776,open_n777,open_n778,open_n779,open_n780,open_n781,open_n782,inst_dob_i16_014}));
  // address_offset=8192;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_008192_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n783,open_n784,open_n785,open_n786,open_n787,open_n788,open_n789,dia[15],open_n790}),
    .dob({open_n815,open_n816,open_n817,open_n818,open_n819,open_n820,open_n821,open_n822,inst_dob_i16_015}));
  // address_offset=9216;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_009216_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i18_008,inst_dob_i18_007,inst_dob_i18_006,inst_dob_i18_005,inst_dob_i18_004,inst_dob_i18_003,inst_dob_i18_002,inst_dob_i18_001,inst_dob_i18_000}));
  // address_offset=10240;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_010240_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i20_008,inst_dob_i20_007,inst_dob_i20_006,inst_dob_i20_005,inst_dob_i20_004,inst_dob_i20_003,inst_dob_i20_002,inst_dob_i20_001,inst_dob_i20_000}));
  // address_offset=11264;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_011264_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i22_008,inst_dob_i22_007,inst_dob_i22_006,inst_dob_i22_005,inst_dob_i22_004,inst_dob_i22_003,inst_dob_i22_002,inst_dob_i22_001,inst_dob_i22_000}));
  // address_offset=12288;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_012288_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i24_008,inst_dob_i24_007,inst_dob_i24_006,inst_dob_i24_005,inst_dob_i24_004,inst_dob_i24_003,inst_dob_i24_002,inst_dob_i24_001,inst_dob_i24_000}));
  // address_offset=13312;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_013312_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i26_008,inst_dob_i26_007,inst_dob_i26_006,inst_dob_i26_005,inst_dob_i26_004,inst_dob_i26_003,inst_dob_i26_002,inst_dob_i26_001,inst_dob_i26_000}));
  // address_offset=14336;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_014336_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i28_008,inst_dob_i28_007,inst_dob_i28_006,inst_dob_i28_005,inst_dob_i28_004,inst_dob_i28_003,inst_dob_i28_002,inst_dob_i28_001,inst_dob_i28_000}));
  // address_offset=15360;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_015360_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i30_008,inst_dob_i30_007,inst_dob_i30_006,inst_dob_i30_005,inst_dob_i30_004,inst_dob_i30_003,inst_dob_i30_002,inst_dob_i30_001,inst_dob_i30_000}));
  // address_offset=16384;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o_al_n54 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o_al_n57 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i32_008,inst_dob_i32_007,inst_dob_i32_006,inst_dob_i32_005,inst_dob_i32_004,inst_dob_i32_003,inst_dob_i32_002,inst_dob_i32_001,inst_dob_i32_000}));
  // address_offset=16384;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1015,open_n1016,open_n1017,open_n1018,open_n1019,open_n1020,open_n1021,dia[9],open_n1022}),
    .dob({open_n1047,open_n1048,open_n1049,open_n1050,open_n1051,open_n1052,open_n1053,open_n1054,inst_dob_i32_009}));
  // address_offset=16384;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1055,open_n1056,open_n1057,open_n1058,open_n1059,open_n1060,open_n1061,dia[10],open_n1062}),
    .dob({open_n1087,open_n1088,open_n1089,open_n1090,open_n1091,open_n1092,open_n1093,open_n1094,inst_dob_i32_010}));
  // address_offset=16384;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1095,open_n1096,open_n1097,open_n1098,open_n1099,open_n1100,open_n1101,dia[11],open_n1102}),
    .dob({open_n1127,open_n1128,open_n1129,open_n1130,open_n1131,open_n1132,open_n1133,open_n1134,inst_dob_i32_011}));
  // address_offset=16384;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1135,open_n1136,open_n1137,open_n1138,open_n1139,open_n1140,open_n1141,dia[12],open_n1142}),
    .dob({open_n1167,open_n1168,open_n1169,open_n1170,open_n1171,open_n1172,open_n1173,open_n1174,inst_dob_i32_012}));
  // address_offset=16384;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1175,open_n1176,open_n1177,open_n1178,open_n1179,open_n1180,open_n1181,dia[13],open_n1182}),
    .dob({open_n1207,open_n1208,open_n1209,open_n1210,open_n1211,open_n1212,open_n1213,open_n1214,inst_dob_i32_013}));
  // address_offset=16384;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1215,open_n1216,open_n1217,open_n1218,open_n1219,open_n1220,open_n1221,dia[14],open_n1222}),
    .dob({open_n1247,open_n1248,open_n1249,open_n1250,open_n1251,open_n1252,open_n1253,open_n1254,inst_dob_i32_014}));
  // address_offset=16384;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_016384_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1255,open_n1256,open_n1257,open_n1258,open_n1259,open_n1260,open_n1261,dia[15],open_n1262}),
    .dob({open_n1287,open_n1288,open_n1289,open_n1290,open_n1291,open_n1292,open_n1293,open_n1294,inst_dob_i32_015}));
  // address_offset=17408;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_017408_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o_al_n54 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o_al_n57 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i34_008,inst_dob_i34_007,inst_dob_i34_006,inst_dob_i34_005,inst_dob_i34_004,inst_dob_i34_003,inst_dob_i34_002,inst_dob_i34_001,inst_dob_i34_000}));
  // address_offset=18432;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_018432_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o_al_n54 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o_al_n57 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i36_008,inst_dob_i36_007,inst_dob_i36_006,inst_dob_i36_005,inst_dob_i36_004,inst_dob_i36_003,inst_dob_i36_002,inst_dob_i36_001,inst_dob_i36_000}));
  // address_offset=19456;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_019456_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_Naddr_o_al_n54 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_Naddr_o_al_n57 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i38_008,inst_dob_i38_007,inst_dob_i38_006,inst_dob_i38_005,inst_dob_i38_004,inst_dob_i38_003,inst_dob_i38_002,inst_dob_i38_001,inst_dob_i38_000}));
  // address_offset=20480;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_020480_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o_al_n70 ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o_al_n73 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i40_008,inst_dob_i40_007,inst_dob_i40_006,inst_dob_i40_005,inst_dob_i40_004,inst_dob_i40_003,inst_dob_i40_002,inst_dob_i40_001,inst_dob_i40_000}));
  // address_offset=21504;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_021504_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o_al_n70 ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o_al_n73 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i42_008,inst_dob_i42_007,inst_dob_i42_006,inst_dob_i42_005,inst_dob_i42_004,inst_dob_i42_003,inst_dob_i42_002,inst_dob_i42_001,inst_dob_i42_000}));
  // address_offset=22528;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_022528_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o_al_n70 ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o_al_n73 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i44_008,inst_dob_i44_007,inst_dob_i44_006,inst_dob_i44_005,inst_dob_i44_004,inst_dob_i44_003,inst_dob_i44_002,inst_dob_i44_001,inst_dob_i44_000}));
  // address_offset=23552;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_023552_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_Naddra_o_al_n70 ,addra[11:10]}),
    .csb({\and_addrb[12]_Naddrb_o_al_n73 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i46_008,inst_dob_i46_007,inst_dob_i46_006,inst_dob_i46_005,inst_dob_i46_004,inst_dob_i46_003,inst_dob_i46_002,inst_dob_i46_001,inst_dob_i46_000}));
  // address_offset=24576;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o_al_n86 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o_al_n89 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i48_008,inst_dob_i48_007,inst_dob_i48_006,inst_dob_i48_005,inst_dob_i48_004,inst_dob_i48_003,inst_dob_i48_002,inst_dob_i48_001,inst_dob_i48_000}));
  // address_offset=24576;data_offset=9;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_009 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1487,open_n1488,open_n1489,open_n1490,open_n1491,open_n1492,open_n1493,dia[9],open_n1494}),
    .dob({open_n1519,open_n1520,open_n1521,open_n1522,open_n1523,open_n1524,open_n1525,open_n1526,inst_dob_i48_009}));
  // address_offset=24576;data_offset=10;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_010 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1527,open_n1528,open_n1529,open_n1530,open_n1531,open_n1532,open_n1533,dia[10],open_n1534}),
    .dob({open_n1559,open_n1560,open_n1561,open_n1562,open_n1563,open_n1564,open_n1565,open_n1566,inst_dob_i48_010}));
  // address_offset=24576;data_offset=11;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_011 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1567,open_n1568,open_n1569,open_n1570,open_n1571,open_n1572,open_n1573,dia[11],open_n1574}),
    .dob({open_n1599,open_n1600,open_n1601,open_n1602,open_n1603,open_n1604,open_n1605,open_n1606,inst_dob_i48_011}));
  // address_offset=24576;data_offset=12;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_012 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1607,open_n1608,open_n1609,open_n1610,open_n1611,open_n1612,open_n1613,dia[12],open_n1614}),
    .dob({open_n1639,open_n1640,open_n1641,open_n1642,open_n1643,open_n1644,open_n1645,open_n1646,inst_dob_i48_012}));
  // address_offset=24576;data_offset=13;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_013 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1647,open_n1648,open_n1649,open_n1650,open_n1651,open_n1652,open_n1653,dia[13],open_n1654}),
    .dob({open_n1679,open_n1680,open_n1681,open_n1682,open_n1683,open_n1684,open_n1685,open_n1686,inst_dob_i48_013}));
  // address_offset=24576;data_offset=14;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_014 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1687,open_n1688,open_n1689,open_n1690,open_n1691,open_n1692,open_n1693,dia[14],open_n1694}),
    .dob({open_n1719,open_n1720,open_n1721,open_n1722,open_n1723,open_n1724,open_n1725,open_n1726,inst_dob_i48_014}));
  // address_offset=24576;data_offset=15;depth=8192;width=1;num_section=1;width_per_section=1;section_size=16;working_depth=8192;working_width=1;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("INV"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("INV"),
    .DATA_WIDTH_A("1"),
    .DATA_WIDTH_B("1"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_024576_015 (
    .addra(addra[12:0]),
    .addrb(addrb[12:0]),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa(addra[15:13]),
    .csb(addrb[15:13]),
    .dia({open_n1727,open_n1728,open_n1729,open_n1730,open_n1731,open_n1732,open_n1733,dia[15],open_n1734}),
    .dob({open_n1759,open_n1760,open_n1761,open_n1762,open_n1763,open_n1764,open_n1765,open_n1766,inst_dob_i48_015}));
  // address_offset=25600;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_025600_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o_al_n86 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o_al_n89 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i50_008,inst_dob_i50_007,inst_dob_i50_006,inst_dob_i50_005,inst_dob_i50_004,inst_dob_i50_003,inst_dob_i50_002,inst_dob_i50_001,inst_dob_i50_000}));
  // address_offset=26624;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_026624_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o_al_n86 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o_al_n89 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i52_008,inst_dob_i52_007,inst_dob_i52_006,inst_dob_i52_005,inst_dob_i52_004,inst_dob_i52_003,inst_dob_i52_002,inst_dob_i52_001,inst_dob_i52_000}));
  // address_offset=27648;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_027648_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[12]_addra_o_al_n86 ,addra[11:10]}),
    .csb({\and_Naddrb[12]_addrb_o_al_n89 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i54_008,inst_dob_i54_007,inst_dob_i54_006,inst_dob_i54_005,inst_dob_i54_004,inst_dob_i54_003,inst_dob_i54_002,inst_dob_i54_001,inst_dob_i54_000}));
  // address_offset=28672;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_028672_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o_al_n102 ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o_al_n105 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i56_008,inst_dob_i56_007,inst_dob_i56_006,inst_dob_i56_005,inst_dob_i56_004,inst_dob_i56_003,inst_dob_i56_002,inst_dob_i56_001,inst_dob_i56_000}));
  // address_offset=29696;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_029696_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o_al_n102 ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o_al_n105 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i58_008,inst_dob_i58_007,inst_dob_i58_006,inst_dob_i58_005,inst_dob_i58_004,inst_dob_i58_003,inst_dob_i58_002,inst_dob_i58_001,inst_dob_i58_000}));
  // address_offset=30720;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("INV"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_030720_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o_al_n102 ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o_al_n105 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i60_008,inst_dob_i60_007,inst_dob_i60_006,inst_dob_i60_005,inst_dob_i60_004,inst_dob_i60_003,inst_dob_i60_002,inst_dob_i60_001,inst_dob_i60_000}));
  // address_offset=31744;data_offset=0;depth=1024;width=9;num_section=1;width_per_section=9;section_size=16;working_depth=1024;working_width=9;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CSA0("SIG"),
    .CSA1("SIG"),
    .CSA2("SIG"),
    .CSB0("SIG"),
    .CSB1("SIG"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("9"),
    .DATA_WIDTH_B("9"),
    .MODE("DP8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_031744_000 (
    .addra({addra[9:0],3'b111}),
    .addrb({addrb[9:0],3'b111}),
    .cea(cea),
    .ceb(ceb),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_addra[12]_addra[_o_al_n102 ,addra[11:10]}),
    .csb({\and_addrb[12]_addrb[_o_al_n105 ,addrb[11:10]}),
    .dia(dia[8:0]),
    .dob({inst_dob_i62_008,inst_dob_i62_007,inst_dob_i62_006,inst_dob_i62_005,inst_dob_i62_004,inst_dob_i62_003,inst_dob_i62_002,inst_dob_i62_001,inst_dob_i62_000}));
  // address_offset=32768;data_offset=0;depth=32;width=16;num_section=1;width_per_section=16;section_size=16;working_depth=512;working_width=18;mode_ecc=0;address_step=1;bytes_in_per_section=1;
  EG_PHY_BRAM #(
    .CEAMUX("1"),
    .CEBMUX("1"),
    .CSA0("INV"),
    .CSA1("INV"),
    .CSA2("SIG"),
    .CSB0("INV"),
    .CSB1("INV"),
    .CSB2("SIG"),
    .DATA_WIDTH_A("18"),
    .DATA_WIDTH_B("18"),
    .MODE("PDPW8K"),
    .OCEAMUX("0"),
    .OCEBMUX("0"),
    .REGMODE_A("NOREG"),
    .REGMODE_B("NOREG"),
    .RESETMODE("SYNC"),
    .RSTAMUX("0"),
    .RSTBMUX("0"),
    .WEAMUX("1"),
    .WEBMUX("0"),
    .WRITEMODE_A("NORMAL"),
    .WRITEMODE_B("NORMAL"))
    inst_32800x16_sub_032768_000 (
    .addra({addra[8:0],4'b1111}),
    .addrb({addrb[8:0],4'b1111}),
    .clka(clka),
    .clkb(clkb),
    .csa({\and_Naddra[11]_Naddr_o_and_cea ,addra[10:9]}),
    .csb({\and_Naddrb[11]_Naddr_o_and_ceb ,addrb[10:9]}),
    .dia(dia[8:0]),
    .dib({open_n1937,open_n1938,dia[15:9]}),
    .doa({inst_dob_i64_008,inst_dob_i64_007,inst_dob_i64_006,inst_dob_i64_005,inst_dob_i64_004,inst_dob_i64_003,inst_dob_i64_002,inst_dob_i64_001,inst_dob_i64_000}),
    .dob({open_n1945,open_n1946,inst_dob_i64_015,inst_dob_i64_014,inst_dob_i64_013,inst_dob_i64_012,inst_dob_i64_011,inst_dob_i64_010,inst_dob_i64_009}));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_0  (
    .i0(inst_dob_i0_000),
    .i1(inst_dob_i2_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_1  (
    .i0(inst_dob_i4_000),
    .i1(inst_dob_i6_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_10  (
    .i0(inst_dob_i40_000),
    .i1(inst_dob_i42_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_10 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_11  (
    .i0(inst_dob_i44_000),
    .i1(inst_dob_i46_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_11 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_12  (
    .i0(inst_dob_i48_000),
    .i1(inst_dob_i50_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_12 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_13  (
    .i0(inst_dob_i52_000),
    .i1(inst_dob_i54_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_13 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_14  (
    .i0(inst_dob_i56_000),
    .i1(inst_dob_i58_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_14 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_15  (
    .i0(inst_dob_i60_000),
    .i1(inst_dob_i62_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_15 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_2  (
    .i0(inst_dob_i8_000),
    .i1(inst_dob_i10_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_3  (
    .i0(inst_dob_i12_000),
    .i1(inst_dob_i14_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_4  (
    .i0(inst_dob_i16_000),
    .i1(inst_dob_i18_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_5  (
    .i0(inst_dob_i20_000),
    .i1(inst_dob_i22_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_6  (
    .i0(inst_dob_i24_000),
    .i1(inst_dob_i26_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_7  (
    .i0(inst_dob_i28_000),
    .i1(inst_dob_i30_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_8  (
    .i0(inst_dob_i32_000),
    .i1(inst_dob_i34_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_8 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_1_9  (
    .i0(inst_dob_i36_000),
    .i1(inst_dob_i38_000),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b0/B1_9 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b0/B1_0 ),
    .i1(\inst_dob_mux_b0/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b0/B1_2 ),
    .i1(\inst_dob_mux_b0/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b0/B1_4 ),
    .i1(\inst_dob_mux_b0/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b0/B1_6 ),
    .i1(\inst_dob_mux_b0/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b0/B1_8 ),
    .i1(\inst_dob_mux_b0/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_4 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b0/B1_10 ),
    .i1(\inst_dob_mux_b0/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_5 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b0/B1_12 ),
    .i1(\inst_dob_mux_b0/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_6 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b0/B1_14 ),
    .i1(\inst_dob_mux_b0/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b0/B2_7 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b0/B2_0 ),
    .i1(\inst_dob_mux_b0/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b0/B2_2 ),
    .i1(\inst_dob_mux_b0/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b0/B2_4 ),
    .i1(\inst_dob_mux_b0/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_2 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b0/B2_6 ),
    .i1(\inst_dob_mux_b0/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b0/B3_3 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b0/B3_0 ),
    .i1(\inst_dob_mux_b0/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b0/B4_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b0/B3_2 ),
    .i1(\inst_dob_mux_b0/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b0/B4_1 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b0/B4_0 ),
    .i1(\inst_dob_mux_b0/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b0/B5_0 ));
  AL_MUX \inst_dob_mux_b0/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b0/B5_0 ),
    .i1(inst_dob_i64_000),
    .sel(addrb_piped[6]),
    .o(dob[0]));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_0  (
    .i0(inst_dob_i0_001),
    .i1(inst_dob_i2_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_1  (
    .i0(inst_dob_i4_001),
    .i1(inst_dob_i6_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_10  (
    .i0(inst_dob_i40_001),
    .i1(inst_dob_i42_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_10 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_11  (
    .i0(inst_dob_i44_001),
    .i1(inst_dob_i46_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_11 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_12  (
    .i0(inst_dob_i48_001),
    .i1(inst_dob_i50_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_12 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_13  (
    .i0(inst_dob_i52_001),
    .i1(inst_dob_i54_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_13 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_14  (
    .i0(inst_dob_i56_001),
    .i1(inst_dob_i58_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_14 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_15  (
    .i0(inst_dob_i60_001),
    .i1(inst_dob_i62_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_15 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_2  (
    .i0(inst_dob_i8_001),
    .i1(inst_dob_i10_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_3  (
    .i0(inst_dob_i12_001),
    .i1(inst_dob_i14_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_4  (
    .i0(inst_dob_i16_001),
    .i1(inst_dob_i18_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_5  (
    .i0(inst_dob_i20_001),
    .i1(inst_dob_i22_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_6  (
    .i0(inst_dob_i24_001),
    .i1(inst_dob_i26_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_7  (
    .i0(inst_dob_i28_001),
    .i1(inst_dob_i30_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_8  (
    .i0(inst_dob_i32_001),
    .i1(inst_dob_i34_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_8 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_1_9  (
    .i0(inst_dob_i36_001),
    .i1(inst_dob_i38_001),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b1/B1_9 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b1/B1_0 ),
    .i1(\inst_dob_mux_b1/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b1/B1_2 ),
    .i1(\inst_dob_mux_b1/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b1/B1_4 ),
    .i1(\inst_dob_mux_b1/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b1/B1_6 ),
    .i1(\inst_dob_mux_b1/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b1/B1_8 ),
    .i1(\inst_dob_mux_b1/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_4 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b1/B1_10 ),
    .i1(\inst_dob_mux_b1/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_5 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b1/B1_12 ),
    .i1(\inst_dob_mux_b1/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_6 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b1/B1_14 ),
    .i1(\inst_dob_mux_b1/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b1/B2_7 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b1/B2_0 ),
    .i1(\inst_dob_mux_b1/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b1/B2_2 ),
    .i1(\inst_dob_mux_b1/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b1/B2_4 ),
    .i1(\inst_dob_mux_b1/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_2 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b1/B2_6 ),
    .i1(\inst_dob_mux_b1/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b1/B3_3 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b1/B3_0 ),
    .i1(\inst_dob_mux_b1/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b1/B4_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b1/B3_2 ),
    .i1(\inst_dob_mux_b1/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b1/B4_1 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b1/B4_0 ),
    .i1(\inst_dob_mux_b1/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b1/B5_0 ));
  AL_MUX \inst_dob_mux_b1/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b1/B5_0 ),
    .i1(inst_dob_i64_001),
    .sel(addrb_piped[6]),
    .o(dob[1]));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_0  (
    .i0(inst_dob_i0_010),
    .i1(inst_dob_i16_010),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b10/B4_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_4_1  (
    .i0(inst_dob_i32_010),
    .i1(inst_dob_i48_010),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b10/B4_1 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b10/B4_0 ),
    .i1(\inst_dob_mux_b10/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b10/B5_0 ));
  AL_MUX \inst_dob_mux_b10/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b10/B5_0 ),
    .i1(inst_dob_i64_010),
    .sel(addrb_piped[6]),
    .o(dob[10]));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_0  (
    .i0(inst_dob_i0_011),
    .i1(inst_dob_i16_011),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b11/B4_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_4_1  (
    .i0(inst_dob_i32_011),
    .i1(inst_dob_i48_011),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b11/B4_1 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b11/B4_0 ),
    .i1(\inst_dob_mux_b11/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b11/B5_0 ));
  AL_MUX \inst_dob_mux_b11/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b11/B5_0 ),
    .i1(inst_dob_i64_011),
    .sel(addrb_piped[6]),
    .o(dob[11]));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_0  (
    .i0(inst_dob_i0_012),
    .i1(inst_dob_i16_012),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b12/B4_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_4_1  (
    .i0(inst_dob_i32_012),
    .i1(inst_dob_i48_012),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b12/B4_1 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b12/B4_0 ),
    .i1(\inst_dob_mux_b12/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b12/B5_0 ));
  AL_MUX \inst_dob_mux_b12/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b12/B5_0 ),
    .i1(inst_dob_i64_012),
    .sel(addrb_piped[6]),
    .o(dob[12]));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_0  (
    .i0(inst_dob_i0_013),
    .i1(inst_dob_i16_013),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b13/B4_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_4_1  (
    .i0(inst_dob_i32_013),
    .i1(inst_dob_i48_013),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b13/B4_1 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b13/B4_0 ),
    .i1(\inst_dob_mux_b13/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b13/B5_0 ));
  AL_MUX \inst_dob_mux_b13/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b13/B5_0 ),
    .i1(inst_dob_i64_013),
    .sel(addrb_piped[6]),
    .o(dob[13]));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_0  (
    .i0(inst_dob_i0_014),
    .i1(inst_dob_i16_014),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b14/B4_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_4_1  (
    .i0(inst_dob_i32_014),
    .i1(inst_dob_i48_014),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b14/B4_1 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b14/B4_0 ),
    .i1(\inst_dob_mux_b14/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b14/B5_0 ));
  AL_MUX \inst_dob_mux_b14/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b14/B5_0 ),
    .i1(inst_dob_i64_014),
    .sel(addrb_piped[6]),
    .o(dob[14]));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_0  (
    .i0(inst_dob_i0_015),
    .i1(inst_dob_i16_015),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b15/B4_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_4_1  (
    .i0(inst_dob_i32_015),
    .i1(inst_dob_i48_015),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b15/B4_1 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b15/B4_0 ),
    .i1(\inst_dob_mux_b15/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b15/B5_0 ));
  AL_MUX \inst_dob_mux_b15/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b15/B5_0 ),
    .i1(inst_dob_i64_015),
    .sel(addrb_piped[6]),
    .o(dob[15]));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_0  (
    .i0(inst_dob_i0_002),
    .i1(inst_dob_i2_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_1  (
    .i0(inst_dob_i4_002),
    .i1(inst_dob_i6_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_10  (
    .i0(inst_dob_i40_002),
    .i1(inst_dob_i42_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_10 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_11  (
    .i0(inst_dob_i44_002),
    .i1(inst_dob_i46_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_11 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_12  (
    .i0(inst_dob_i48_002),
    .i1(inst_dob_i50_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_12 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_13  (
    .i0(inst_dob_i52_002),
    .i1(inst_dob_i54_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_13 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_14  (
    .i0(inst_dob_i56_002),
    .i1(inst_dob_i58_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_14 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_15  (
    .i0(inst_dob_i60_002),
    .i1(inst_dob_i62_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_15 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_2  (
    .i0(inst_dob_i8_002),
    .i1(inst_dob_i10_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_3  (
    .i0(inst_dob_i12_002),
    .i1(inst_dob_i14_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_4  (
    .i0(inst_dob_i16_002),
    .i1(inst_dob_i18_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_5  (
    .i0(inst_dob_i20_002),
    .i1(inst_dob_i22_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_6  (
    .i0(inst_dob_i24_002),
    .i1(inst_dob_i26_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_7  (
    .i0(inst_dob_i28_002),
    .i1(inst_dob_i30_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_8  (
    .i0(inst_dob_i32_002),
    .i1(inst_dob_i34_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_8 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_1_9  (
    .i0(inst_dob_i36_002),
    .i1(inst_dob_i38_002),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b2/B1_9 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b2/B1_0 ),
    .i1(\inst_dob_mux_b2/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b2/B1_2 ),
    .i1(\inst_dob_mux_b2/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b2/B1_4 ),
    .i1(\inst_dob_mux_b2/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b2/B1_6 ),
    .i1(\inst_dob_mux_b2/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b2/B1_8 ),
    .i1(\inst_dob_mux_b2/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_4 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b2/B1_10 ),
    .i1(\inst_dob_mux_b2/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_5 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b2/B1_12 ),
    .i1(\inst_dob_mux_b2/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_6 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b2/B1_14 ),
    .i1(\inst_dob_mux_b2/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b2/B2_7 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b2/B2_0 ),
    .i1(\inst_dob_mux_b2/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b2/B2_2 ),
    .i1(\inst_dob_mux_b2/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b2/B2_4 ),
    .i1(\inst_dob_mux_b2/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_2 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b2/B2_6 ),
    .i1(\inst_dob_mux_b2/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b2/B3_3 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b2/B3_0 ),
    .i1(\inst_dob_mux_b2/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b2/B4_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b2/B3_2 ),
    .i1(\inst_dob_mux_b2/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b2/B4_1 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b2/B4_0 ),
    .i1(\inst_dob_mux_b2/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b2/B5_0 ));
  AL_MUX \inst_dob_mux_b2/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b2/B5_0 ),
    .i1(inst_dob_i64_002),
    .sel(addrb_piped[6]),
    .o(dob[2]));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_0  (
    .i0(inst_dob_i0_003),
    .i1(inst_dob_i2_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_1  (
    .i0(inst_dob_i4_003),
    .i1(inst_dob_i6_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_10  (
    .i0(inst_dob_i40_003),
    .i1(inst_dob_i42_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_10 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_11  (
    .i0(inst_dob_i44_003),
    .i1(inst_dob_i46_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_11 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_12  (
    .i0(inst_dob_i48_003),
    .i1(inst_dob_i50_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_12 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_13  (
    .i0(inst_dob_i52_003),
    .i1(inst_dob_i54_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_13 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_14  (
    .i0(inst_dob_i56_003),
    .i1(inst_dob_i58_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_14 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_15  (
    .i0(inst_dob_i60_003),
    .i1(inst_dob_i62_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_15 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_2  (
    .i0(inst_dob_i8_003),
    .i1(inst_dob_i10_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_3  (
    .i0(inst_dob_i12_003),
    .i1(inst_dob_i14_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_4  (
    .i0(inst_dob_i16_003),
    .i1(inst_dob_i18_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_5  (
    .i0(inst_dob_i20_003),
    .i1(inst_dob_i22_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_6  (
    .i0(inst_dob_i24_003),
    .i1(inst_dob_i26_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_7  (
    .i0(inst_dob_i28_003),
    .i1(inst_dob_i30_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_8  (
    .i0(inst_dob_i32_003),
    .i1(inst_dob_i34_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_8 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_1_9  (
    .i0(inst_dob_i36_003),
    .i1(inst_dob_i38_003),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b3/B1_9 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b3/B1_0 ),
    .i1(\inst_dob_mux_b3/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b3/B1_2 ),
    .i1(\inst_dob_mux_b3/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b3/B1_4 ),
    .i1(\inst_dob_mux_b3/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b3/B1_6 ),
    .i1(\inst_dob_mux_b3/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b3/B1_8 ),
    .i1(\inst_dob_mux_b3/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_4 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b3/B1_10 ),
    .i1(\inst_dob_mux_b3/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_5 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b3/B1_12 ),
    .i1(\inst_dob_mux_b3/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_6 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b3/B1_14 ),
    .i1(\inst_dob_mux_b3/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b3/B2_7 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b3/B2_0 ),
    .i1(\inst_dob_mux_b3/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b3/B2_2 ),
    .i1(\inst_dob_mux_b3/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b3/B2_4 ),
    .i1(\inst_dob_mux_b3/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_2 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b3/B2_6 ),
    .i1(\inst_dob_mux_b3/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b3/B3_3 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b3/B3_0 ),
    .i1(\inst_dob_mux_b3/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b3/B4_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b3/B3_2 ),
    .i1(\inst_dob_mux_b3/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b3/B4_1 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b3/B4_0 ),
    .i1(\inst_dob_mux_b3/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b3/B5_0 ));
  AL_MUX \inst_dob_mux_b3/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b3/B5_0 ),
    .i1(inst_dob_i64_003),
    .sel(addrb_piped[6]),
    .o(dob[3]));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_0  (
    .i0(inst_dob_i0_004),
    .i1(inst_dob_i2_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_1  (
    .i0(inst_dob_i4_004),
    .i1(inst_dob_i6_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_10  (
    .i0(inst_dob_i40_004),
    .i1(inst_dob_i42_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_10 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_11  (
    .i0(inst_dob_i44_004),
    .i1(inst_dob_i46_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_11 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_12  (
    .i0(inst_dob_i48_004),
    .i1(inst_dob_i50_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_12 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_13  (
    .i0(inst_dob_i52_004),
    .i1(inst_dob_i54_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_13 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_14  (
    .i0(inst_dob_i56_004),
    .i1(inst_dob_i58_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_14 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_15  (
    .i0(inst_dob_i60_004),
    .i1(inst_dob_i62_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_15 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_2  (
    .i0(inst_dob_i8_004),
    .i1(inst_dob_i10_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_3  (
    .i0(inst_dob_i12_004),
    .i1(inst_dob_i14_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_4  (
    .i0(inst_dob_i16_004),
    .i1(inst_dob_i18_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_5  (
    .i0(inst_dob_i20_004),
    .i1(inst_dob_i22_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_6  (
    .i0(inst_dob_i24_004),
    .i1(inst_dob_i26_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_7  (
    .i0(inst_dob_i28_004),
    .i1(inst_dob_i30_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_8  (
    .i0(inst_dob_i32_004),
    .i1(inst_dob_i34_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_8 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_1_9  (
    .i0(inst_dob_i36_004),
    .i1(inst_dob_i38_004),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b4/B1_9 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b4/B1_0 ),
    .i1(\inst_dob_mux_b4/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b4/B1_2 ),
    .i1(\inst_dob_mux_b4/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b4/B1_4 ),
    .i1(\inst_dob_mux_b4/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b4/B1_6 ),
    .i1(\inst_dob_mux_b4/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b4/B1_8 ),
    .i1(\inst_dob_mux_b4/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_4 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b4/B1_10 ),
    .i1(\inst_dob_mux_b4/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_5 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b4/B1_12 ),
    .i1(\inst_dob_mux_b4/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_6 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b4/B1_14 ),
    .i1(\inst_dob_mux_b4/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b4/B2_7 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b4/B2_0 ),
    .i1(\inst_dob_mux_b4/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b4/B2_2 ),
    .i1(\inst_dob_mux_b4/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b4/B2_4 ),
    .i1(\inst_dob_mux_b4/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_2 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b4/B2_6 ),
    .i1(\inst_dob_mux_b4/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b4/B3_3 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b4/B3_0 ),
    .i1(\inst_dob_mux_b4/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b4/B4_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b4/B3_2 ),
    .i1(\inst_dob_mux_b4/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b4/B4_1 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b4/B4_0 ),
    .i1(\inst_dob_mux_b4/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b4/B5_0 ));
  AL_MUX \inst_dob_mux_b4/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b4/B5_0 ),
    .i1(inst_dob_i64_004),
    .sel(addrb_piped[6]),
    .o(dob[4]));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_0  (
    .i0(inst_dob_i0_005),
    .i1(inst_dob_i2_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_1  (
    .i0(inst_dob_i4_005),
    .i1(inst_dob_i6_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_10  (
    .i0(inst_dob_i40_005),
    .i1(inst_dob_i42_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_10 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_11  (
    .i0(inst_dob_i44_005),
    .i1(inst_dob_i46_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_11 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_12  (
    .i0(inst_dob_i48_005),
    .i1(inst_dob_i50_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_12 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_13  (
    .i0(inst_dob_i52_005),
    .i1(inst_dob_i54_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_13 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_14  (
    .i0(inst_dob_i56_005),
    .i1(inst_dob_i58_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_14 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_15  (
    .i0(inst_dob_i60_005),
    .i1(inst_dob_i62_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_15 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_2  (
    .i0(inst_dob_i8_005),
    .i1(inst_dob_i10_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_3  (
    .i0(inst_dob_i12_005),
    .i1(inst_dob_i14_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_4  (
    .i0(inst_dob_i16_005),
    .i1(inst_dob_i18_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_5  (
    .i0(inst_dob_i20_005),
    .i1(inst_dob_i22_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_6  (
    .i0(inst_dob_i24_005),
    .i1(inst_dob_i26_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_7  (
    .i0(inst_dob_i28_005),
    .i1(inst_dob_i30_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_8  (
    .i0(inst_dob_i32_005),
    .i1(inst_dob_i34_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_8 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_1_9  (
    .i0(inst_dob_i36_005),
    .i1(inst_dob_i38_005),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b5/B1_9 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b5/B1_0 ),
    .i1(\inst_dob_mux_b5/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b5/B1_2 ),
    .i1(\inst_dob_mux_b5/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b5/B1_4 ),
    .i1(\inst_dob_mux_b5/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b5/B1_6 ),
    .i1(\inst_dob_mux_b5/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b5/B1_8 ),
    .i1(\inst_dob_mux_b5/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_4 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b5/B1_10 ),
    .i1(\inst_dob_mux_b5/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_5 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b5/B1_12 ),
    .i1(\inst_dob_mux_b5/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_6 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b5/B1_14 ),
    .i1(\inst_dob_mux_b5/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b5/B2_7 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b5/B2_0 ),
    .i1(\inst_dob_mux_b5/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b5/B2_2 ),
    .i1(\inst_dob_mux_b5/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b5/B2_4 ),
    .i1(\inst_dob_mux_b5/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_2 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b5/B2_6 ),
    .i1(\inst_dob_mux_b5/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b5/B3_3 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b5/B3_0 ),
    .i1(\inst_dob_mux_b5/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b5/B4_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b5/B3_2 ),
    .i1(\inst_dob_mux_b5/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b5/B4_1 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b5/B4_0 ),
    .i1(\inst_dob_mux_b5/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b5/B5_0 ));
  AL_MUX \inst_dob_mux_b5/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b5/B5_0 ),
    .i1(inst_dob_i64_005),
    .sel(addrb_piped[6]),
    .o(dob[5]));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_0  (
    .i0(inst_dob_i0_006),
    .i1(inst_dob_i2_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_1  (
    .i0(inst_dob_i4_006),
    .i1(inst_dob_i6_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_10  (
    .i0(inst_dob_i40_006),
    .i1(inst_dob_i42_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_10 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_11  (
    .i0(inst_dob_i44_006),
    .i1(inst_dob_i46_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_11 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_12  (
    .i0(inst_dob_i48_006),
    .i1(inst_dob_i50_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_12 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_13  (
    .i0(inst_dob_i52_006),
    .i1(inst_dob_i54_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_13 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_14  (
    .i0(inst_dob_i56_006),
    .i1(inst_dob_i58_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_14 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_15  (
    .i0(inst_dob_i60_006),
    .i1(inst_dob_i62_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_15 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_2  (
    .i0(inst_dob_i8_006),
    .i1(inst_dob_i10_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_3  (
    .i0(inst_dob_i12_006),
    .i1(inst_dob_i14_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_4  (
    .i0(inst_dob_i16_006),
    .i1(inst_dob_i18_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_5  (
    .i0(inst_dob_i20_006),
    .i1(inst_dob_i22_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_6  (
    .i0(inst_dob_i24_006),
    .i1(inst_dob_i26_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_7  (
    .i0(inst_dob_i28_006),
    .i1(inst_dob_i30_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_8  (
    .i0(inst_dob_i32_006),
    .i1(inst_dob_i34_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_8 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_1_9  (
    .i0(inst_dob_i36_006),
    .i1(inst_dob_i38_006),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b6/B1_9 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b6/B1_0 ),
    .i1(\inst_dob_mux_b6/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b6/B1_2 ),
    .i1(\inst_dob_mux_b6/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b6/B1_4 ),
    .i1(\inst_dob_mux_b6/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b6/B1_6 ),
    .i1(\inst_dob_mux_b6/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b6/B1_8 ),
    .i1(\inst_dob_mux_b6/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_4 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b6/B1_10 ),
    .i1(\inst_dob_mux_b6/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_5 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b6/B1_12 ),
    .i1(\inst_dob_mux_b6/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_6 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b6/B1_14 ),
    .i1(\inst_dob_mux_b6/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b6/B2_7 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b6/B2_0 ),
    .i1(\inst_dob_mux_b6/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b6/B2_2 ),
    .i1(\inst_dob_mux_b6/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b6/B2_4 ),
    .i1(\inst_dob_mux_b6/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_2 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b6/B2_6 ),
    .i1(\inst_dob_mux_b6/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b6/B3_3 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b6/B3_0 ),
    .i1(\inst_dob_mux_b6/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b6/B4_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b6/B3_2 ),
    .i1(\inst_dob_mux_b6/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b6/B4_1 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b6/B4_0 ),
    .i1(\inst_dob_mux_b6/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b6/B5_0 ));
  AL_MUX \inst_dob_mux_b6/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b6/B5_0 ),
    .i1(inst_dob_i64_006),
    .sel(addrb_piped[6]),
    .o(dob[6]));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_0  (
    .i0(inst_dob_i0_007),
    .i1(inst_dob_i2_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_1  (
    .i0(inst_dob_i4_007),
    .i1(inst_dob_i6_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_10  (
    .i0(inst_dob_i40_007),
    .i1(inst_dob_i42_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_10 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_11  (
    .i0(inst_dob_i44_007),
    .i1(inst_dob_i46_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_11 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_12  (
    .i0(inst_dob_i48_007),
    .i1(inst_dob_i50_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_12 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_13  (
    .i0(inst_dob_i52_007),
    .i1(inst_dob_i54_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_13 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_14  (
    .i0(inst_dob_i56_007),
    .i1(inst_dob_i58_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_14 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_15  (
    .i0(inst_dob_i60_007),
    .i1(inst_dob_i62_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_15 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_2  (
    .i0(inst_dob_i8_007),
    .i1(inst_dob_i10_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_3  (
    .i0(inst_dob_i12_007),
    .i1(inst_dob_i14_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_4  (
    .i0(inst_dob_i16_007),
    .i1(inst_dob_i18_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_5  (
    .i0(inst_dob_i20_007),
    .i1(inst_dob_i22_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_6  (
    .i0(inst_dob_i24_007),
    .i1(inst_dob_i26_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_7  (
    .i0(inst_dob_i28_007),
    .i1(inst_dob_i30_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_8  (
    .i0(inst_dob_i32_007),
    .i1(inst_dob_i34_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_8 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_1_9  (
    .i0(inst_dob_i36_007),
    .i1(inst_dob_i38_007),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b7/B1_9 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b7/B1_0 ),
    .i1(\inst_dob_mux_b7/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b7/B1_2 ),
    .i1(\inst_dob_mux_b7/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b7/B1_4 ),
    .i1(\inst_dob_mux_b7/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b7/B1_6 ),
    .i1(\inst_dob_mux_b7/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b7/B1_8 ),
    .i1(\inst_dob_mux_b7/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_4 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b7/B1_10 ),
    .i1(\inst_dob_mux_b7/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_5 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b7/B1_12 ),
    .i1(\inst_dob_mux_b7/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_6 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b7/B1_14 ),
    .i1(\inst_dob_mux_b7/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b7/B2_7 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b7/B2_0 ),
    .i1(\inst_dob_mux_b7/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b7/B2_2 ),
    .i1(\inst_dob_mux_b7/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b7/B2_4 ),
    .i1(\inst_dob_mux_b7/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_2 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b7/B2_6 ),
    .i1(\inst_dob_mux_b7/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b7/B3_3 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b7/B3_0 ),
    .i1(\inst_dob_mux_b7/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b7/B4_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b7/B3_2 ),
    .i1(\inst_dob_mux_b7/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b7/B4_1 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b7/B4_0 ),
    .i1(\inst_dob_mux_b7/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b7/B5_0 ));
  AL_MUX \inst_dob_mux_b7/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b7/B5_0 ),
    .i1(inst_dob_i64_007),
    .sel(addrb_piped[6]),
    .o(dob[7]));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_0  (
    .i0(inst_dob_i0_008),
    .i1(inst_dob_i2_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_1  (
    .i0(inst_dob_i4_008),
    .i1(inst_dob_i6_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_10  (
    .i0(inst_dob_i40_008),
    .i1(inst_dob_i42_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_10 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_11  (
    .i0(inst_dob_i44_008),
    .i1(inst_dob_i46_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_11 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_12  (
    .i0(inst_dob_i48_008),
    .i1(inst_dob_i50_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_12 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_13  (
    .i0(inst_dob_i52_008),
    .i1(inst_dob_i54_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_13 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_14  (
    .i0(inst_dob_i56_008),
    .i1(inst_dob_i58_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_14 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_15  (
    .i0(inst_dob_i60_008),
    .i1(inst_dob_i62_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_15 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_2  (
    .i0(inst_dob_i8_008),
    .i1(inst_dob_i10_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_3  (
    .i0(inst_dob_i12_008),
    .i1(inst_dob_i14_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_4  (
    .i0(inst_dob_i16_008),
    .i1(inst_dob_i18_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_5  (
    .i0(inst_dob_i20_008),
    .i1(inst_dob_i22_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_6  (
    .i0(inst_dob_i24_008),
    .i1(inst_dob_i26_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_7  (
    .i0(inst_dob_i28_008),
    .i1(inst_dob_i30_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_8  (
    .i0(inst_dob_i32_008),
    .i1(inst_dob_i34_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_8 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_1_9  (
    .i0(inst_dob_i36_008),
    .i1(inst_dob_i38_008),
    .sel(addrb_piped[1]),
    .o(\inst_dob_mux_b8/B1_9 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_0  (
    .i0(\inst_dob_mux_b8/B1_0 ),
    .i1(\inst_dob_mux_b8/B1_1 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_1  (
    .i0(\inst_dob_mux_b8/B1_2 ),
    .i1(\inst_dob_mux_b8/B1_3 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_2  (
    .i0(\inst_dob_mux_b8/B1_4 ),
    .i1(\inst_dob_mux_b8/B1_5 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_3  (
    .i0(\inst_dob_mux_b8/B1_6 ),
    .i1(\inst_dob_mux_b8/B1_7 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_4  (
    .i0(\inst_dob_mux_b8/B1_8 ),
    .i1(\inst_dob_mux_b8/B1_9 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_4 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_5  (
    .i0(\inst_dob_mux_b8/B1_10 ),
    .i1(\inst_dob_mux_b8/B1_11 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_5 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_6  (
    .i0(\inst_dob_mux_b8/B1_12 ),
    .i1(\inst_dob_mux_b8/B1_13 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_6 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_2_7  (
    .i0(\inst_dob_mux_b8/B1_14 ),
    .i1(\inst_dob_mux_b8/B1_15 ),
    .sel(addrb_piped[2]),
    .o(\inst_dob_mux_b8/B2_7 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_0  (
    .i0(\inst_dob_mux_b8/B2_0 ),
    .i1(\inst_dob_mux_b8/B2_1 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_1  (
    .i0(\inst_dob_mux_b8/B2_2 ),
    .i1(\inst_dob_mux_b8/B2_3 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_2  (
    .i0(\inst_dob_mux_b8/B2_4 ),
    .i1(\inst_dob_mux_b8/B2_5 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_2 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_3_3  (
    .i0(\inst_dob_mux_b8/B2_6 ),
    .i1(\inst_dob_mux_b8/B2_7 ),
    .sel(addrb_piped[3]),
    .o(\inst_dob_mux_b8/B3_3 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_0  (
    .i0(\inst_dob_mux_b8/B3_0 ),
    .i1(\inst_dob_mux_b8/B3_1 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b8/B4_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_4_1  (
    .i0(\inst_dob_mux_b8/B3_2 ),
    .i1(\inst_dob_mux_b8/B3_3 ),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b8/B4_1 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b8/B4_0 ),
    .i1(\inst_dob_mux_b8/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b8/B5_0 ));
  AL_MUX \inst_dob_mux_b8/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b8/B5_0 ),
    .i1(inst_dob_i64_008),
    .sel(addrb_piped[6]),
    .o(dob[8]));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_0  (
    .i0(inst_dob_i0_009),
    .i1(inst_dob_i16_009),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b9/B4_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_4_1  (
    .i0(inst_dob_i32_009),
    .i1(inst_dob_i48_009),
    .sel(addrb_piped[4]),
    .o(\inst_dob_mux_b9/B4_1 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_5_0  (
    .i0(\inst_dob_mux_b9/B4_0 ),
    .i1(\inst_dob_mux_b9/B4_1 ),
    .sel(addrb_piped[5]),
    .o(\inst_dob_mux_b9/B5_0 ));
  AL_MUX \inst_dob_mux_b9/al_mux_b0_6_0  (
    .i0(\inst_dob_mux_b9/B5_0 ),
    .i1(inst_dob_i64_009),
    .sel(addrb_piped[6]),
    .o(dob[9]));

endmodule 

module AL_DFF_X
  (
  ar,
  as,
  clk,
  d,
  en,
  sr,
  ss,
  q
  );

  input ar;
  input as;
  input clk;
  input d;
  input en;
  input sr;
  input ss;
  output q;

  wire enout;
  wire srout;
  wire ssout;

  AL_MUX u_en (
    .i0(q),
    .i1(d),
    .sel(en),
    .o(enout));
  AL_MUX u_reset (
    .i0(ssout),
    .i1(1'b0),
    .sel(sr),
    .o(srout));
  AL_DFF u_seq (
    .clk(clk),
    .d(srout),
    .reset(ar),
    .set(as),
    .q(q));
  AL_MUX u_set (
    .i0(enout),
    .i1(1'b1),
    .sel(ss),
    .o(ssout));

endmodule 

module AL_MUX
  (
  input i0,
  input i1,
  input sel,
  output o
  );

  wire not_sel, sel_i0, sel_i1;
  not u0 (not_sel, sel);
  and u1 (sel_i1, sel, i1);
  and u2 (sel_i0, not_sel, i0);
  or u3 (o, sel_i1, sel_i0);

endmodule

module AL_DFF
  (
  input reset,
  input set,
  input clk,
  input d,
  output reg q
  );

  parameter INI = 1'b0;

  // synthesis translate_off
  tri0 gsrn = glbl.gsrn;

  always @(gsrn)
  begin
    if(!gsrn)
      assign q = INI;
    else
      deassign q;
  end
  // synthesis translate_on

  always @(posedge reset or posedge set or posedge clk)
  begin
    if (reset)
      q <= 1'b0;
    else if (set)
      q <= 1'b1;
    else
      q <= d;
  end

endmodule

